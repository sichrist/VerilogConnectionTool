

module testmodule_a
(

	input in1,
	input in2,
	output out

	);

	endmodule