

module testmodule_b
(


	input in1,
	input in2,
	output out

	);

	testmodule_c testinstance
	(

	);

	endmodule