module testmodule_c(

	input in1,
	input in2,
	output out

	);


	endmodule
